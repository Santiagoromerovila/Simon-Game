library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package trabajo_pkg is
 
  type std_logic_array is array (0 to 7) of std_logic_vector(1 downto 0);
  
end package trabajo_pkg;
 
-- Package Body Section
package body trabajo_pkg is

end package body trabajo_pkg;